// File: Arch.bsv
package Arch;
typedef 64 DATA_WIDTH;
Integer data_width = valueOf(DATA_WIDTH);
endpackage
